module final(LED, INPUT);
	input INPUT;
	output LED;
	assign LED = INPUT;
	
endmodule
